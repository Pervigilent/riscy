parameter FIFO_PTR_CHIPYZ_CHANNEL0    = 5,
          FIFO_WIDTH_CHIPXYZ_CHANNEL0 = 32;

parameter FIFO_PTR_CHIPYZ_CHANNEL1    = 6,
          FIFO_WIDTH_CHIPXYZ_CHANNEL1 = 32;

parameter FIFO_PTR_CHIPYZ_CHANNEL2    = 8,
          FIFO_WIDTH_CHIPXYZ_CHANNEL2 = 16;
