module rcv_c (
	rcv_c_in1,
	rcv_c_in2,
	rcv_c_in3,
	rcv_c_out1,
	rcv_c_out2
);
	// --------------------
	input rcv_c_in1;
	input [7:0] rcv_c_in2;
	input rcv_c_in3;
	output [7:0] rcv_c_out1;
	output rcv_c_out2;
	// --------------------
	// Synthesizable RTL code
	always @(*) begin
		// -----
		// -----
	end
end module

