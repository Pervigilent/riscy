module rcv_d (
    rcv_d_in1,
    rcv_d_in2,
    rcv_d_out1,
    rcv_d_out2,
    rcv_d_in3
);
    // --------------------
    input        rcv_d_in1;
    input        rcv_d_in2;

    output       rcv_d_out1;
    output [7:0] rcv_d_out2;
    output       rcv_d_out3;
    // --------------------
    // Synthesizable RTL code
    always @(*) begin
        // -----
        // -----
    end
end module

