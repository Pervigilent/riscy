module xmit_b (
	xmit_b_in1,
	xmit_b_in2,
	xmit_b_in3,
	xmit_b_out1,
	xmit_b_out2
);
	// --------------------
	input [7:0] xmit_b_in1;
	input xmit_b_in2;
	input xmit_b_in3;
	output xmit_b_out1;
	output xmit_b_out2;
	// --------------------
	// Synthesizable RTL code
	always @(*) begin
		// -----
		// -----
	end
end module

